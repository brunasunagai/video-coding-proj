library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.type_pack.all;

entity cl_sad_8x8_parallel is 
port(
    ori: in input_64;
    ref: in input_64;
    sad_out: out std_logic_vector(14 downto 0)
);
end cl_sad_8x8_parallel;

architecture arch_sad of cl_sad_8x8_parallel is 

-- Components 
component adder is 
 generic (N: integer);
 port(
 		A, B: in std_logic_vector(N-1 downto 0);
 		S: out std_logic_vector(N downto 0)
 );
 end component; 


-- Signals
signal neg_ref_0: std_logic_vector(7 downto 0);
signal neg_ref_1: std_logic_vector(7 downto 0);
signal neg_ref_2: std_logic_vector(7 downto 0);
signal neg_ref_3: std_logic_vector(7 downto 0);
signal neg_ref_4: std_logic_vector(7 downto 0);
signal neg_ref_5: std_logic_vector(7 downto 0);
signal neg_ref_6: std_logic_vector(7 downto 0);
signal neg_ref_7: std_logic_vector(7 downto 0);
signal neg_ref_8: std_logic_vector(7 downto 0);
signal neg_ref_9: std_logic_vector(7 downto 0);
signal neg_ref_10: std_logic_vector(7 downto 0);
signal neg_ref_11: std_logic_vector(7 downto 0);
signal neg_ref_12: std_logic_vector(7 downto 0);
signal neg_ref_13: std_logic_vector(7 downto 0);
signal neg_ref_14: std_logic_vector(7 downto 0);
signal neg_ref_15: std_logic_vector(7 downto 0);
signal neg_ref_16: std_logic_vector(7 downto 0);
signal neg_ref_17: std_logic_vector(7 downto 0);
signal neg_ref_18: std_logic_vector(7 downto 0);
signal neg_ref_19: std_logic_vector(7 downto 0);
signal neg_ref_20: std_logic_vector(7 downto 0);
signal neg_ref_21: std_logic_vector(7 downto 0);
signal neg_ref_22: std_logic_vector(7 downto 0);
signal neg_ref_23: std_logic_vector(7 downto 0);
signal neg_ref_24: std_logic_vector(7 downto 0);
signal neg_ref_25: std_logic_vector(7 downto 0);
signal neg_ref_26: std_logic_vector(7 downto 0);
signal neg_ref_27: std_logic_vector(7 downto 0);
signal neg_ref_28: std_logic_vector(7 downto 0);
signal neg_ref_29: std_logic_vector(7 downto 0);
signal neg_ref_30: std_logic_vector(7 downto 0);
signal neg_ref_31: std_logic_vector(7 downto 0);
signal neg_ref_32: std_logic_vector(7 downto 0);
signal neg_ref_33: std_logic_vector(7 downto 0);
signal neg_ref_34: std_logic_vector(7 downto 0);
signal neg_ref_35: std_logic_vector(7 downto 0);
signal neg_ref_36: std_logic_vector(7 downto 0);
signal neg_ref_37: std_logic_vector(7 downto 0);
signal neg_ref_38: std_logic_vector(7 downto 0);
signal neg_ref_39: std_logic_vector(7 downto 0);
signal neg_ref_40: std_logic_vector(7 downto 0);
signal neg_ref_41: std_logic_vector(7 downto 0);
signal neg_ref_42: std_logic_vector(7 downto 0);
signal neg_ref_43: std_logic_vector(7 downto 0);
signal neg_ref_44: std_logic_vector(7 downto 0);
signal neg_ref_45: std_logic_vector(7 downto 0);
signal neg_ref_46: std_logic_vector(7 downto 0);
signal neg_ref_47: std_logic_vector(7 downto 0);
signal neg_ref_48: std_logic_vector(7 downto 0);
signal neg_ref_49: std_logic_vector(7 downto 0);
signal neg_ref_50: std_logic_vector(7 downto 0);
signal neg_ref_51: std_logic_vector(7 downto 0);
signal neg_ref_52: std_logic_vector(7 downto 0);
signal neg_ref_53: std_logic_vector(7 downto 0);
signal neg_ref_54: std_logic_vector(7 downto 0);
signal neg_ref_55: std_logic_vector(7 downto 0);
signal neg_ref_56: std_logic_vector(7 downto 0);
signal neg_ref_57: std_logic_vector(7 downto 0);
signal neg_ref_58: std_logic_vector(7 downto 0);
signal neg_ref_59: std_logic_vector(7 downto 0);
signal neg_ref_60: std_logic_vector(7 downto 0);
signal neg_ref_61: std_logic_vector(7 downto 0);
signal neg_ref_62: std_logic_vector(7 downto 0);
signal neg_ref_63: std_logic_vector(7 downto 0);

signal sub_0: std_logic_vector(8 downto 0);
signal sub_1: std_logic_vector(8 downto 0);
signal sub_2: std_logic_vector(8 downto 0);
signal sub_3: std_logic_vector(8 downto 0);
signal sub_4: std_logic_vector(8 downto 0);
signal sub_5: std_logic_vector(8 downto 0);
signal sub_6: std_logic_vector(8 downto 0);
signal sub_7: std_logic_vector(8 downto 0);
signal sub_8: std_logic_vector(8 downto 0);
signal sub_9: std_logic_vector(8 downto 0);
signal sub_10: std_logic_vector(8 downto 0);
signal sub_11: std_logic_vector(8 downto 0);
signal sub_12: std_logic_vector(8 downto 0);
signal sub_13: std_logic_vector(8 downto 0);
signal sub_14: std_logic_vector(8 downto 0);
signal sub_15: std_logic_vector(8 downto 0);
signal sub_16: std_logic_vector(8 downto 0);
signal sub_17: std_logic_vector(8 downto 0);
signal sub_18: std_logic_vector(8 downto 0);
signal sub_19: std_logic_vector(8 downto 0);
signal sub_20: std_logic_vector(8 downto 0);
signal sub_21: std_logic_vector(8 downto 0);
signal sub_22: std_logic_vector(8 downto 0);
signal sub_23: std_logic_vector(8 downto 0);
signal sub_24: std_logic_vector(8 downto 0);
signal sub_25: std_logic_vector(8 downto 0);
signal sub_26: std_logic_vector(8 downto 0);
signal sub_27: std_logic_vector(8 downto 0);
signal sub_28: std_logic_vector(8 downto 0);
signal sub_29: std_logic_vector(8 downto 0);
signal sub_30: std_logic_vector(8 downto 0);
signal sub_31: std_logic_vector(8 downto 0);
signal sub_32: std_logic_vector(8 downto 0);
signal sub_33: std_logic_vector(8 downto 0);
signal sub_34: std_logic_vector(8 downto 0);
signal sub_35: std_logic_vector(8 downto 0);
signal sub_36: std_logic_vector(8 downto 0);
signal sub_37: std_logic_vector(8 downto 0);
signal sub_38: std_logic_vector(8 downto 0);
signal sub_39: std_logic_vector(8 downto 0);
signal sub_40: std_logic_vector(8 downto 0);
signal sub_41: std_logic_vector(8 downto 0);
signal sub_42: std_logic_vector(8 downto 0);
signal sub_43: std_logic_vector(8 downto 0);
signal sub_44: std_logic_vector(8 downto 0);
signal sub_45: std_logic_vector(8 downto 0);
signal sub_46: std_logic_vector(8 downto 0);
signal sub_47: std_logic_vector(8 downto 0);
signal sub_48: std_logic_vector(8 downto 0);
signal sub_49: std_logic_vector(8 downto 0);
signal sub_50: std_logic_vector(8 downto 0);
signal sub_51: std_logic_vector(8 downto 0);
signal sub_52: std_logic_vector(8 downto 0);
signal sub_53: std_logic_vector(8 downto 0);
signal sub_54: std_logic_vector(8 downto 0);
signal sub_55: std_logic_vector(8 downto 0);
signal sub_56: std_logic_vector(8 downto 0);
signal sub_57: std_logic_vector(8 downto 0);
signal sub_58: std_logic_vector(8 downto 0);
signal sub_59: std_logic_vector(8 downto 0);
signal sub_60: std_logic_vector(8 downto 0);
signal sub_61: std_logic_vector(8 downto 0);
signal sub_62: std_logic_vector(8 downto 0);
signal sub_63: std_logic_vector(8 downto 0);

signal abs_0: std_logic_vector(8 downto 0);
signal abs_1: std_logic_vector(8 downto 0);
signal abs_2: std_logic_vector(8 downto 0);
signal abs_3: std_logic_vector(8 downto 0);
signal abs_4: std_logic_vector(8 downto 0);
signal abs_5: std_logic_vector(8 downto 0);
signal abs_6: std_logic_vector(8 downto 0);
signal abs_7: std_logic_vector(8 downto 0);
signal abs_8: std_logic_vector(8 downto 0);
signal abs_9: std_logic_vector(8 downto 0);
signal abs_10: std_logic_vector(8 downto 0);
signal abs_11: std_logic_vector(8 downto 0);
signal abs_12: std_logic_vector(8 downto 0);
signal abs_13: std_logic_vector(8 downto 0);
signal abs_14: std_logic_vector(8 downto 0);
signal abs_15: std_logic_vector(8 downto 0);
signal abs_16: std_logic_vector(8 downto 0);
signal abs_17: std_logic_vector(8 downto 0);
signal abs_18: std_logic_vector(8 downto 0);
signal abs_19: std_logic_vector(8 downto 0);
signal abs_20: std_logic_vector(8 downto 0);
signal abs_21: std_logic_vector(8 downto 0);
signal abs_22: std_logic_vector(8 downto 0);
signal abs_23: std_logic_vector(8 downto 0);
signal abs_24: std_logic_vector(8 downto 0);
signal abs_25: std_logic_vector(8 downto 0);
signal abs_26: std_logic_vector(8 downto 0);
signal abs_27: std_logic_vector(8 downto 0);
signal abs_28: std_logic_vector(8 downto 0);
signal abs_29: std_logic_vector(8 downto 0);
signal abs_30: std_logic_vector(8 downto 0);
signal abs_31: std_logic_vector(8 downto 0);
signal abs_32: std_logic_vector(8 downto 0);
signal abs_33: std_logic_vector(8 downto 0);
signal abs_34: std_logic_vector(8 downto 0);
signal abs_35: std_logic_vector(8 downto 0);
signal abs_36: std_logic_vector(8 downto 0);
signal abs_37: std_logic_vector(8 downto 0);
signal abs_38: std_logic_vector(8 downto 0);
signal abs_39: std_logic_vector(8 downto 0);
signal abs_40: std_logic_vector(8 downto 0);
signal abs_41: std_logic_vector(8 downto 0);
signal abs_42: std_logic_vector(8 downto 0);
signal abs_43: std_logic_vector(8 downto 0);
signal abs_44: std_logic_vector(8 downto 0);
signal abs_45: std_logic_vector(8 downto 0);
signal abs_46: std_logic_vector(8 downto 0);
signal abs_47: std_logic_vector(8 downto 0);
signal abs_48: std_logic_vector(8 downto 0);
signal abs_49: std_logic_vector(8 downto 0);
signal abs_50: std_logic_vector(8 downto 0);
signal abs_51: std_logic_vector(8 downto 0);
signal abs_52: std_logic_vector(8 downto 0);
signal abs_53: std_logic_vector(8 downto 0);
signal abs_54: std_logic_vector(8 downto 0);
signal abs_55: std_logic_vector(8 downto 0);
signal abs_56: std_logic_vector(8 downto 0);
signal abs_57: std_logic_vector(8 downto 0);
signal abs_58: std_logic_vector(8 downto 0);
signal abs_59: std_logic_vector(8 downto 0);
signal abs_60: std_logic_vector(8 downto 0);
signal abs_61: std_logic_vector(8 downto 0);
signal abs_62: std_logic_vector(8 downto 0);
signal abs_63: std_logic_vector(8 downto 0);

signal sum_01: std_logic_vector(9 downto 0);
signal sum_23: std_logic_vector(9 downto 0);
signal sum_45: std_logic_vector(9 downto 0);
signal sum_67: std_logic_vector(9 downto 0);
signal sum_89: std_logic_vector(9 downto 0);
signal sum_1011: std_logic_vector(9 downto 0);
signal sum_1213: std_logic_vector(9 downto 0);
signal sum_1415: std_logic_vector(9 downto 0);
signal sum_1617: std_logic_vector(9 downto 0);
signal sum_1819: std_logic_vector(9 downto 0);
signal sum_2021: std_logic_vector(9 downto 0);
signal sum_2223: std_logic_vector(9 downto 0);
signal sum_2425: std_logic_vector(9 downto 0);
signal sum_2627: std_logic_vector(9 downto 0);
signal sum_2829: std_logic_vector(9 downto 0);
signal sum_3031: std_logic_vector(9 downto 0);
signal sum_3233: std_logic_vector(9 downto 0);
signal sum_3435: std_logic_vector(9 downto 0);
signal sum_3637: std_logic_vector(9 downto 0);
signal sum_3839: std_logic_vector(9 downto 0);
signal sum_4041: std_logic_vector(9 downto 0);
signal sum_4243: std_logic_vector(9 downto 0);
signal sum_4445: std_logic_vector(9 downto 0);
signal sum_4647: std_logic_vector(9 downto 0);
signal sum_4849: std_logic_vector(9 downto 0);
signal sum_5051: std_logic_vector(9 downto 0);
signal sum_5253: std_logic_vector(9 downto 0);
signal sum_5455: std_logic_vector(9 downto 0);
signal sum_5657: std_logic_vector(9 downto 0);
signal sum_5859: std_logic_vector(9 downto 0);
signal sum_6061: std_logic_vector(9 downto 0);
signal sum_6263: std_logic_vector(9 downto 0);

signal sum_after_10: std_logic_vector(10 downto 0);
signal sum_after_11: std_logic_vector(10 downto 0);
signal sum_after_12: std_logic_vector(10 downto 0);
signal sum_after_13: std_logic_vector(10 downto 0);
signal sum_after_14: std_logic_vector(10 downto 0);
signal sum_after_15: std_logic_vector(10 downto 0);
signal sum_after_16: std_logic_vector(10 downto 0);
signal sum_after_17: std_logic_vector(10 downto 0);
signal sum_after_18: std_logic_vector(10 downto 0);
signal sum_after_19: std_logic_vector(10 downto 0);
signal sum_after_110: std_logic_vector(10 downto 0);
signal sum_after_111: std_logic_vector(10 downto 0);
signal sum_after_112: std_logic_vector(10 downto 0);
signal sum_after_113: std_logic_vector(10 downto 0);
signal sum_after_114: std_logic_vector(10 downto 0);
signal sum_after_115: std_logic_vector(10 downto 0);
signal sum_after_20: std_logic_vector(11 downto 0);
signal sum_after_21: std_logic_vector(11 downto 0);
signal sum_after_22: std_logic_vector(11 downto 0);
signal sum_after_23: std_logic_vector(11 downto 0);
signal sum_after_24: std_logic_vector(11 downto 0);
signal sum_after_25: std_logic_vector(11 downto 0);
signal sum_after_26: std_logic_vector(11 downto 0);
signal sum_after_27: std_logic_vector(11 downto 0);
signal sum_after_30: std_logic_vector(12 downto 0);
signal sum_after_31: std_logic_vector(12 downto 0);
signal sum_after_32: std_logic_vector(12 downto 0);
signal sum_after_33: std_logic_vector(12 downto 0);
signal sum_after_40: std_logic_vector(13 downto 0);
signal sum_after_41: std_logic_vector(13 downto 0);
signal sum_after_50: std_logic_vector(14 downto 0);


begin

neg_ref_0 <= std_logic_vector(resize(-signed(ref(0)),8));
neg_ref_1 <= std_logic_vector(resize(-signed(ref(1)),8));
neg_ref_2 <= std_logic_vector(resize(-signed(ref(2)),8));
neg_ref_3 <= std_logic_vector(resize(-signed(ref(3)),8));
neg_ref_4 <= std_logic_vector(resize(-signed(ref(4)),8));
neg_ref_5 <= std_logic_vector(resize(-signed(ref(5)),8));
neg_ref_6 <= std_logic_vector(resize(-signed(ref(6)),8));
neg_ref_7 <= std_logic_vector(resize(-signed(ref(7)),8));
neg_ref_8 <= std_logic_vector(resize(-signed(ref(8)),8));
neg_ref_9 <= std_logic_vector(resize(-signed(ref(9)),8));
neg_ref_10 <= std_logic_vector(resize(-signed(ref(10)),8));
neg_ref_11 <= std_logic_vector(resize(-signed(ref(11)),8));
neg_ref_12 <= std_logic_vector(resize(-signed(ref(12)),8));
neg_ref_13 <= std_logic_vector(resize(-signed(ref(13)),8));
neg_ref_14 <= std_logic_vector(resize(-signed(ref(14)),8));
neg_ref_15 <= std_logic_vector(resize(-signed(ref(15)),8));
neg_ref_16 <= std_logic_vector(resize(-signed(ref(16)),8));
neg_ref_17 <= std_logic_vector(resize(-signed(ref(17)),8));
neg_ref_18 <= std_logic_vector(resize(-signed(ref(18)),8));
neg_ref_19 <= std_logic_vector(resize(-signed(ref(19)),8));
neg_ref_20 <= std_logic_vector(resize(-signed(ref(20)),8));
neg_ref_21 <= std_logic_vector(resize(-signed(ref(21)),8));
neg_ref_22 <= std_logic_vector(resize(-signed(ref(22)),8));
neg_ref_23 <= std_logic_vector(resize(-signed(ref(23)),8));
neg_ref_24 <= std_logic_vector(resize(-signed(ref(24)),8));
neg_ref_25 <= std_logic_vector(resize(-signed(ref(25)),8));
neg_ref_26 <= std_logic_vector(resize(-signed(ref(26)),8));
neg_ref_27 <= std_logic_vector(resize(-signed(ref(27)),8));
neg_ref_28 <= std_logic_vector(resize(-signed(ref(28)),8));
neg_ref_29 <= std_logic_vector(resize(-signed(ref(29)),8));
neg_ref_30 <= std_logic_vector(resize(-signed(ref(30)),8));
neg_ref_31 <= std_logic_vector(resize(-signed(ref(31)),8));
neg_ref_32 <= std_logic_vector(resize(-signed(ref(32)),8));
neg_ref_33 <= std_logic_vector(resize(-signed(ref(33)),8));
neg_ref_34 <= std_logic_vector(resize(-signed(ref(34)),8));
neg_ref_35 <= std_logic_vector(resize(-signed(ref(35)),8));
neg_ref_36 <= std_logic_vector(resize(-signed(ref(36)),8));
neg_ref_37 <= std_logic_vector(resize(-signed(ref(37)),8));
neg_ref_38 <= std_logic_vector(resize(-signed(ref(38)),8));
neg_ref_39 <= std_logic_vector(resize(-signed(ref(39)),8));
neg_ref_40 <= std_logic_vector(resize(-signed(ref(40)),8));
neg_ref_41 <= std_logic_vector(resize(-signed(ref(41)),8));
neg_ref_42 <= std_logic_vector(resize(-signed(ref(42)),8));
neg_ref_43 <= std_logic_vector(resize(-signed(ref(43)),8));
neg_ref_44 <= std_logic_vector(resize(-signed(ref(44)),8));
neg_ref_45 <= std_logic_vector(resize(-signed(ref(45)),8));
neg_ref_46 <= std_logic_vector(resize(-signed(ref(46)),8));
neg_ref_47 <= std_logic_vector(resize(-signed(ref(47)),8));
neg_ref_48 <= std_logic_vector(resize(-signed(ref(48)),8));
neg_ref_49 <= std_logic_vector(resize(-signed(ref(49)),8));
neg_ref_50 <= std_logic_vector(resize(-signed(ref(50)),8));
neg_ref_51 <= std_logic_vector(resize(-signed(ref(51)),8));
neg_ref_52 <= std_logic_vector(resize(-signed(ref(52)),8));
neg_ref_53 <= std_logic_vector(resize(-signed(ref(53)),8));
neg_ref_54 <= std_logic_vector(resize(-signed(ref(54)),8));
neg_ref_55 <= std_logic_vector(resize(-signed(ref(55)),8));
neg_ref_56 <= std_logic_vector(resize(-signed(ref(56)),8));
neg_ref_57 <= std_logic_vector(resize(-signed(ref(57)),8));
neg_ref_58 <= std_logic_vector(resize(-signed(ref(58)),8));
neg_ref_59 <= std_logic_vector(resize(-signed(ref(59)),8));
neg_ref_60 <= std_logic_vector(resize(-signed(ref(60)),8));
neg_ref_61 <= std_logic_vector(resize(-signed(ref(61)),8));
neg_ref_62 <= std_logic_vector(resize(-signed(ref(62)),8));
neg_ref_63 <= std_logic_vector(resize(-signed(ref(63)),8));

abs_0 <= std_logic_vector(abs(signed(sub_0)));
abs_1 <= std_logic_vector(abs(signed(sub_1)));
abs_2 <= std_logic_vector(abs(signed(sub_2)));
abs_3 <= std_logic_vector(abs(signed(sub_3)));
abs_4 <= std_logic_vector(abs(signed(sub_4)));
abs_5 <= std_logic_vector(abs(signed(sub_5)));
abs_6 <= std_logic_vector(abs(signed(sub_6)));
abs_7 <= std_logic_vector(abs(signed(sub_7)));
abs_8 <= std_logic_vector(abs(signed(sub_8)));
abs_9 <= std_logic_vector(abs(signed(sub_9)));
abs_10 <= std_logic_vector(abs(signed(sub_10)));
abs_11 <= std_logic_vector(abs(signed(sub_11)));
abs_12 <= std_logic_vector(abs(signed(sub_12)));
abs_13 <= std_logic_vector(abs(signed(sub_13)));
abs_14 <= std_logic_vector(abs(signed(sub_14)));
abs_15 <= std_logic_vector(abs(signed(sub_15)));
abs_16 <= std_logic_vector(abs(signed(sub_16)));
abs_17 <= std_logic_vector(abs(signed(sub_17)));
abs_18 <= std_logic_vector(abs(signed(sub_18)));
abs_19 <= std_logic_vector(abs(signed(sub_19)));
abs_20 <= std_logic_vector(abs(signed(sub_20)));
abs_21 <= std_logic_vector(abs(signed(sub_21)));
abs_22 <= std_logic_vector(abs(signed(sub_22)));
abs_23 <= std_logic_vector(abs(signed(sub_23)));
abs_24 <= std_logic_vector(abs(signed(sub_24)));
abs_25 <= std_logic_vector(abs(signed(sub_25)));
abs_26 <= std_logic_vector(abs(signed(sub_26)));
abs_27 <= std_logic_vector(abs(signed(sub_27)));
abs_28 <= std_logic_vector(abs(signed(sub_28)));
abs_29 <= std_logic_vector(abs(signed(sub_29)));
abs_30 <= std_logic_vector(abs(signed(sub_30)));
abs_31 <= std_logic_vector(abs(signed(sub_31)));
abs_32 <= std_logic_vector(abs(signed(sub_32)));
abs_33 <= std_logic_vector(abs(signed(sub_33)));
abs_34 <= std_logic_vector(abs(signed(sub_34)));
abs_35 <= std_logic_vector(abs(signed(sub_35)));
abs_36 <= std_logic_vector(abs(signed(sub_36)));
abs_37 <= std_logic_vector(abs(signed(sub_37)));
abs_38 <= std_logic_vector(abs(signed(sub_38)));
abs_39 <= std_logic_vector(abs(signed(sub_39)));
abs_40 <= std_logic_vector(abs(signed(sub_40)));
abs_41 <= std_logic_vector(abs(signed(sub_41)));
abs_42 <= std_logic_vector(abs(signed(sub_42)));
abs_43 <= std_logic_vector(abs(signed(sub_43)));
abs_44 <= std_logic_vector(abs(signed(sub_44)));
abs_45 <= std_logic_vector(abs(signed(sub_45)));
abs_46 <= std_logic_vector(abs(signed(sub_46)));
abs_47 <= std_logic_vector(abs(signed(sub_47)));
abs_48 <= std_logic_vector(abs(signed(sub_48)));
abs_49 <= std_logic_vector(abs(signed(sub_49)));
abs_50 <= std_logic_vector(abs(signed(sub_50)));
abs_51 <= std_logic_vector(abs(signed(sub_51)));
abs_52 <= std_logic_vector(abs(signed(sub_52)));
abs_53 <= std_logic_vector(abs(signed(sub_53)));
abs_54 <= std_logic_vector(abs(signed(sub_54)));
abs_55 <= std_logic_vector(abs(signed(sub_55)));
abs_56 <= std_logic_vector(abs(signed(sub_56)));
abs_57 <= std_logic_vector(abs(signed(sub_57)));
abs_58 <= std_logic_vector(abs(signed(sub_58)));
abs_59 <= std_logic_vector(abs(signed(sub_59)));
abs_60 <= std_logic_vector(abs(signed(sub_60)));
abs_61 <= std_logic_vector(abs(signed(sub_61)));
abs_62 <= std_logic_vector(abs(signed(sub_62)));
abs_63 <= std_logic_vector(abs(signed(sub_63)));


SUB0: adder generic map (8) port map (ori(0),neg_ref_0,sub_0);
SUB1: adder generic map (8) port map (ori(1),neg_ref_1,sub_1);
SUB2: adder generic map (8) port map (ori(2),neg_ref_2,sub_2);
SUB3: adder generic map (8) port map (ori(3),neg_ref_3,sub_3);
SUB4: adder generic map (8) port map (ori(4),neg_ref_4,sub_4);
SUB5: adder generic map (8) port map (ori(5),neg_ref_5,sub_5);
SUB6: adder generic map (8) port map (ori(6),neg_ref_6,sub_6);
SUB7: adder generic map (8) port map (ori(7),neg_ref_7,sub_7);
SUB8: adder generic map (8) port map (ori(8),neg_ref_8,sub_8);
SUB9: adder generic map (8) port map (ori(9),neg_ref_9,sub_9);
SUB10: adder generic map (8) port map (ori(10),neg_ref_10,sub_10);
SUB11: adder generic map (8) port map (ori(11),neg_ref_11,sub_11);
SUB12: adder generic map (8) port map (ori(12),neg_ref_12,sub_12);
SUB13: adder generic map (8) port map (ori(13),neg_ref_13,sub_13);
SUB14: adder generic map (8) port map (ori(14),neg_ref_14,sub_14);
SUB15: adder generic map (8) port map (ori(15),neg_ref_15,sub_15);
SUB16: adder generic map (8) port map (ori(16),neg_ref_16,sub_16);
SUB17: adder generic map (8) port map (ori(17),neg_ref_17,sub_17);
SUB18: adder generic map (8) port map (ori(18),neg_ref_18,sub_18);
SUB19: adder generic map (8) port map (ori(19),neg_ref_19,sub_19);
SUB20: adder generic map (8) port map (ori(20),neg_ref_20,sub_20);
SUB21: adder generic map (8) port map (ori(21),neg_ref_21,sub_21);
SUB22: adder generic map (8) port map (ori(22),neg_ref_22,sub_22);
SUB23: adder generic map (8) port map (ori(23),neg_ref_23,sub_23);
SUB24: adder generic map (8) port map (ori(24),neg_ref_24,sub_24);
SUB25: adder generic map (8) port map (ori(25),neg_ref_25,sub_25);
SUB26: adder generic map (8) port map (ori(26),neg_ref_26,sub_26);
SUB27: adder generic map (8) port map (ori(27),neg_ref_27,sub_27);
SUB28: adder generic map (8) port map (ori(28),neg_ref_28,sub_28);
SUB29: adder generic map (8) port map (ori(29),neg_ref_29,sub_29);
SUB30: adder generic map (8) port map (ori(30),neg_ref_30,sub_30);
SUB31: adder generic map (8) port map (ori(31),neg_ref_31,sub_31);
SUB32: adder generic map (8) port map (ori(32),neg_ref_32,sub_32);
SUB33: adder generic map (8) port map (ori(33),neg_ref_33,sub_33);
SUB34: adder generic map (8) port map (ori(34),neg_ref_34,sub_34);
SUB35: adder generic map (8) port map (ori(35),neg_ref_35,sub_35);
SUB36: adder generic map (8) port map (ori(36),neg_ref_36,sub_36);
SUB37: adder generic map (8) port map (ori(37),neg_ref_37,sub_37);
SUB38: adder generic map (8) port map (ori(38),neg_ref_38,sub_38);
SUB39: adder generic map (8) port map (ori(39),neg_ref_39,sub_39);
SUB40: adder generic map (8) port map (ori(40),neg_ref_40,sub_40);
SUB41: adder generic map (8) port map (ori(41),neg_ref_41,sub_41);
SUB42: adder generic map (8) port map (ori(42),neg_ref_42,sub_42);
SUB43: adder generic map (8) port map (ori(43),neg_ref_43,sub_43);
SUB44: adder generic map (8) port map (ori(44),neg_ref_44,sub_44);
SUB45: adder generic map (8) port map (ori(45),neg_ref_45,sub_45);
SUB46: adder generic map (8) port map (ori(46),neg_ref_46,sub_46);
SUB47: adder generic map (8) port map (ori(47),neg_ref_47,sub_47);
SUB48: adder generic map (8) port map (ori(48),neg_ref_48,sub_48);
SUB49: adder generic map (8) port map (ori(49),neg_ref_49,sub_49);
SUB50: adder generic map (8) port map (ori(50),neg_ref_50,sub_50);
SUB51: adder generic map (8) port map (ori(51),neg_ref_51,sub_51);
SUB52: adder generic map (8) port map (ori(52),neg_ref_52,sub_52);
SUB53: adder generic map (8) port map (ori(53),neg_ref_53,sub_53);
SUB54: adder generic map (8) port map (ori(54),neg_ref_54,sub_54);
SUB55: adder generic map (8) port map (ori(55),neg_ref_55,sub_55);
SUB56: adder generic map (8) port map (ori(56),neg_ref_56,sub_56);
SUB57: adder generic map (8) port map (ori(57),neg_ref_57,sub_57);
SUB58: adder generic map (8) port map (ori(58),neg_ref_58,sub_58);
SUB59: adder generic map (8) port map (ori(59),neg_ref_59,sub_59);
SUB60: adder generic map (8) port map (ori(60),neg_ref_60,sub_60);
SUB61: adder generic map (8) port map (ori(61),neg_ref_61,sub_61);
SUB62: adder generic map (8) port map (ori(62),neg_ref_62,sub_62);
SUB63: adder generic map (8) port map (ori(63),neg_ref_63,sub_63);

ADD00: adder generic map (9) port map (abs_0,abs_1,sum_01);
ADD01: adder generic map (9) port map (abs_2,abs_3,sum_23);
ADD02: adder generic map (9) port map (abs_4,abs_5,sum_45);
ADD03: adder generic map (9) port map (abs_6,abs_7,sum_67);
ADD04: adder generic map (9) port map (abs_8,abs_9,sum_89);
ADD05: adder generic map (9) port map (abs_10,abs_11,sum_1011);
ADD06: adder generic map (9) port map (abs_12,abs_13,sum_1213);
ADD07: adder generic map (9) port map (abs_14,abs_15,sum_1415);
ADD08: adder generic map (9) port map (abs_16,abs_17,sum_1617);
ADD09: adder generic map (9) port map (abs_18,abs_19,sum_1819);
ADD010: adder generic map (9) port map (abs_20,abs_21,sum_2021);
ADD011: adder generic map (9) port map (abs_22,abs_23,sum_2223);
ADD012: adder generic map (9) port map (abs_24,abs_25,sum_2425);
ADD013: adder generic map (9) port map (abs_26,abs_27,sum_2627);
ADD014: adder generic map (9) port map (abs_28,abs_29,sum_2829);
ADD015: adder generic map (9) port map (abs_30,abs_31,sum_3031);
ADD016: adder generic map (9) port map (abs_32,abs_33,sum_3233);
ADD017: adder generic map (9) port map (abs_34,abs_35,sum_3435);
ADD018: adder generic map (9) port map (abs_36,abs_37,sum_3637);
ADD019: adder generic map (9) port map (abs_38,abs_39,sum_3839);
ADD020: adder generic map (9) port map (abs_40,abs_41,sum_4041);
ADD021: adder generic map (9) port map (abs_42,abs_43,sum_4243);
ADD022: adder generic map (9) port map (abs_44,abs_45,sum_4445);
ADD023: adder generic map (9) port map (abs_46,abs_47,sum_4647);
ADD024: adder generic map (9) port map (abs_48,abs_49,sum_4849);
ADD025: adder generic map (9) port map (abs_50,abs_51,sum_5051);
ADD026: adder generic map (9) port map (abs_52,abs_53,sum_5253);
ADD027: adder generic map (9) port map (abs_54,abs_55,sum_5455);
ADD028: adder generic map (9) port map (abs_56,abs_57,sum_5657);
ADD029: adder generic map (9) port map (abs_58,abs_59,sum_5859);
ADD030: adder generic map (9) port map (abs_60,abs_61,sum_6061);
ADD031: adder generic map (9) port map (abs_62,abs_63,sum_6263);

ADD10: adder generic map (10) port map (sum_01,sum_23,sum_after_10);
ADD11: adder generic map (10) port map (sum_45,sum_67,sum_after_11);
ADD12: adder generic map (10) port map (sum_89,sum_1011,sum_after_12);
ADD13: adder generic map (10) port map (sum_1213,sum_1415,sum_after_13);
ADD14: adder generic map (10) port map (sum_1617,sum_1819,sum_after_14);
ADD15: adder generic map (10) port map (sum_2021,sum_2223,sum_after_15);
ADD16: adder generic map (10) port map (sum_2425,sum_2627,sum_after_16);
ADD17: adder generic map (10) port map (sum_2829,sum_3031,sum_after_17);
ADD18: adder generic map (10) port map (sum_3233,sum_3435,sum_after_18);
ADD19: adder generic map (10) port map (sum_3637,sum_3839,sum_after_19);
ADD110: adder generic map (10) port map (sum_4041,sum_4243,sum_after_110);
ADD111: adder generic map (10) port map (sum_4445,sum_4647,sum_after_111);
ADD112: adder generic map (10) port map (sum_4849,sum_5051,sum_after_112);
ADD113: adder generic map (10) port map (sum_5253,sum_5455,sum_after_113);
ADD114: adder generic map (10) port map (sum_5657,sum_5859,sum_after_114);
ADD115: adder generic map (10) port map (sum_6061,sum_6263,sum_after_115);
ADD20: adder generic map (11) port map (sum_after_10,sum_after_11,sum_after_20);
ADD21: adder generic map (11) port map (sum_after_12,sum_after_13,sum_after_21);
ADD22: adder generic map (11) port map (sum_after_14,sum_after_15,sum_after_22);
ADD23: adder generic map (11) port map (sum_after_16,sum_after_17,sum_after_23);
ADD24: adder generic map (11) port map (sum_after_18,sum_after_19,sum_after_24);
ADD25: adder generic map (11) port map (sum_after_110,sum_after_111,sum_after_25);
ADD26: adder generic map (11) port map (sum_after_112,sum_after_113,sum_after_26);
ADD27: adder generic map (11) port map (sum_after_114,sum_after_115,sum_after_27);
ADD30: adder generic map (12) port map (sum_after_20,sum_after_21,sum_after_30);
ADD31: adder generic map (12) port map (sum_after_22,sum_after_23,sum_after_31);
ADD32: adder generic map (12) port map (sum_after_24,sum_after_25,sum_after_32);
ADD33: adder generic map (12) port map (sum_after_26,sum_after_27,sum_after_33);
ADD40: adder generic map (13) port map (sum_after_30,sum_after_31,sum_after_40);
ADD41: adder generic map (13) port map (sum_after_32,sum_after_33,sum_after_41);
ADD50: adder generic map (14) port map (sum_after_40,sum_after_41,sum_after_50);


sad_out <= sum_after_50;

end arch_sad;